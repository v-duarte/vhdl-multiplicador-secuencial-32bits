library verilog;
use verilog.vl_types.all;
entity MULTIPLICADORSECUENCIAL_vlg_vec_tst is
end MULTIPLICADORSECUENCIAL_vlg_vec_tst;
